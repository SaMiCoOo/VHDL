library IEEE;
use IEEE.std_logic_1164.all;

entity write_decoder is
	port(
		i:	in std_logic_vector(3 downto 0);
		o0,o1,o2,o3,
		o4,o5,o6,o7,
		o8,o9,o10,o11,
		o12,o13,o14,o15:	out std_logic
	);
end write_decoder;

architecture behavior of write_decoder is
begin
 	process(i)
	begin
		case i is
			when "0000"=> 
		o0<= '1';	o1<= '0';	o2<= '0';	o3<= '0';
		o4<= '0';	o5<= '0';	o6<= '0';	o7<= '0';
		o8<= '0';	o9<= '0';	o10<= '0';	o11<= '0';
		o12<= '0';	o13<= '0';	o14<= '0';	o15<= '0';
			when "0001"=> 
		o0<= '0';	o1<= '1';	o2<= '0';	o3<= '0';
		o4<= '0';	o5<= '0';	o6<= '0';	o7<= '0';
		o8<= '0';	o9<= '0';	o10<= '0';	o11<= '0';
		o12<= '0';	o13<= '0';	o14<= '0';	o15<= '0';
			when "0010"=> 
		o0<= '0';	o1<= '0';	o2<= '1';	o3<= '0';
		o4<= '0';	o5<= '0';	o6<= '0';	o7<= '0';
		o8<= '0';	o9<= '0';	o10<= '0';	o11<= '0';
		o12<= '0';	o13<= '0';	o14<= '0';	o15<= '0';
			when "0011"=> 
		o0<= '0';	o1<= '0';	o2<= '0';	o3<= '1';
		o4<= '0';	o5<= '0';	o6<= '0';	o7<= '0';
		o8<= '0';	o9<= '0';	o10<= '0';	o11<= '0';
		o12<= '0';	o13<= '0';	o14<= '0';	o15<= '0';
			when "0100"=> 
		o0<= '0';	o1<= '0';	o2<= '0';	o3<= '0';
		o4<= '1';	o5<= '0';	o6<= '0';	o7<= '0';
		o8<= '0';	o9<= '0';	o10<= '0';	o11<= '0';
		o12<= '0';	o13<= '0';	o14<= '0';	o15<= '0';
			when "0101"=> 
		o0<= '0';	o1<= '0';	o2<= '0';	o3<= '0';
		o4<= '0';	o5<= '1';	o6<= '0';	o7<= '0';
		o8<= '0';	o9<= '0';	o10<= '0';	o11<= '0';
		o12<= '0';	o13<= '0';	o14<= '0';	o15<= '0';
			when "0110"=> 
		o0<= '0';	o1<= '0';	o2<= '0';	o3<= '0';
		o4<= '0';	o5<= '0';	o6<= '1';	o7<= '0';
		o8<= '0';	o9<= '0';	o10<= '0';	o11<= '0';
		o12<= '0';	o13<= '0';	o14<= '0';	o15<= '0';
			when "0111"=> 
		o0<= '0';	o1<= '0';	o2<= '0';	o3<= '0';
		o4<= '0';	o5<= '0';	o6<= '0';	o7<= '1';
		o8<= '0';	o9<= '0';	o10<= '0';	o11<= '0';
		o12<= '0';	o13<= '0';	o14<= '0';	o15<= '0';
			when "1000"=> 
		o0<= '0';	o1<= '0';	o2<= '0';	o3<= '0';
		o4<= '0';	o5<= '0';	o6<= '0';	o7<= '0';
		o8<= '1';	o9<= '0';	o10<= '0';	o11<= '0';
		o12<= '0';	o13<= '0';	o14<= '0';	o15<= '0';
			when "1001"=> 
		o0<= '0';	o1<= '0';	o2<= '0';	o3<= '0';
		o4<= '0';	o5<= '0';	o6<= '0';	o7<= '0';
		o8<= '0';	o9<= '1';	o10<= '0';	o11<= '0';
		o12<= '0';	o13<= '0';	o14<= '0';	o15<= '0';
			when "1010"=> 
		o0<= '0';	o1<= '0';	o2<= '0';	o3<= '0';
		o4<= '0';	o5<= '0';	o6<= '0';	o7<= '0';
		o8<= '0';	o9<= '0';	o10<= '1';	o11<= '0';
		o12<= '0';	o13<= '0';	o14<= '0';	o15<= '0';
			when "1011"=> 
		o0<= '0';	o1<= '0';	o2<= '0';	o3<= '0';
		o4<= '0';	o5<= '0';	o6<= '0';	o7<= '0';
		o8<= '0';	o9<= '0';	o10<= '0';	o11<= '1';
		o12<= '0';	o13<= '0';	o14<= '0';	o15<= '0';
			when "1100"=> 
		o0<= '0';	o1<= '0';	o2<= '0';	o3<= '0';
		o4<= '0';	o5<= '0';	o6<= '0';	o7<= '0';
		o8<= '0';	o9<= '0';	o10<= '0';	o11<= '0';
		o12<= '1';	o13<= '0';	o14<= '0';	o15<= '0';
			when "1101"=> 
		o0<= '0';	o1<= '0';	o2<= '0';	o3<= '0';
		o4<= '0';	o5<= '0';	o6<= '0';	o7<= '0';
		o8<= '0';	o9<= '0';	o10<= '0';	o11<= '0';
		o12<= '0';	o13<= '1';	o14<= '0';	o15<= '0';
			when "1110"=> 
		o0<= '0';	o1<= '0';	o2<= '0';	o3<= '0';
		o4<= '0';	o5<= '0';	o6<= '0';	o7<= '0';
		o8<= '0';	o9<= '0';	o10<= '0';	o11<= '0';
		o12<= '0';	o13<= '0';	o14<= '1';	o15<= '0';
			when "1111"=> 
		o0<= '0';	o1<= '0';	o2<= '0';	o3<= '0';
		o4<= '0';	o5<= '0';	o6<= '0';	o7<= '0';
		o8<= '0';	o9<= '0';	o10<= '0';	o11<= '0';
		o12<= '0';	o13<= '0';	o14<= '0';	o15<= '1';
			when others =>
		o0<= '0';	o1<= '0';	o2<= '0';	o3<= '0';
		o4<= '0';	o5<= '0';	o6<= '0';	o7<= '0';
		o8<= '0';	o9<= '0';	o10<= '0';	o11<= '0';
		o12<= '0';	o13<= '0';	o14<= '0';	o15<= '0';

		end case;
	end process ;
	



end;
